-- VHDL model created from schematic KAZKAS.sch -- Apr 24 17:27:14 2022

library IEEE;
use IEEE.std_logic_1164.all;
library xp2;
use xp2.components.all;

entity KAZKAS is
end KAZKAS;

architecture SCHEMATIC of KAZKAS is

   SIGNAL gnd : std_logic := '0';
   SIGNAL vcc : std_logic := '1';


begin


end SCHEMATIC;
