------------------------------------- 

--KTU 2015

--Informatikos fakultetas
--Kompiuteriu katedra
--Kompiuteriu Architektura [P175B125] 
--Kazimieras Bagdonas 

--v1.0

------------------------------------- 
--KTU 2016 

--ditto

--v1.01
--panaikinta "save" mikrokomanda registrams, sutrumpinta ROM eilute nuo 75 iki 69 bitu, nesuderinama su V1.0   

------------------------------------- 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is 
	port (
		RST_ROM 	: in std_logic;
		clk 		: in std_logic;
		ROM_CMD 	: in std_logic_vector(7 downto 0);  
		ROM_Dout 	: out std_logic_vector(1 to 69)
		);
end ROM ;

architecture rtl of ROM is
	
	type memory is array (0 to 255) of std_logic_vector(1 to 69) ; 
	
	constant ROM_CMDln : memory := (  
--                    1         2         3         4         5         6            Dvi komentaro eilutes duoda bitu numerius   
--           123456789012345678901234567890123456789012345678901234567890123456789    (nuo 1 iki 69)
0=> "010000000000000100000000000000000000000000000000000000000000000000000",  --Komentaro vieta
1=> "010000000000000000000010000001000000000000000000000000000000000000000",  --Komentaro vieta
2=> "010000000000000000000000000000000000100000000000000000000000000000000",  --Komentaro vieta
3=> "000010000000000000000000000000000000000000000000000000000000000000000",  --Komentaro vieta
4=> "110000000011000000000000000000000000000000000000000000000000000000000",  --Komentaro vieta
5=> "000000001000000000000000000000000000000000000000001000000000000000000",  --Komentaro vieta
6=> "000000000000000000000000000000000000000000000000000000000000000000001",  --Komentaro vieta
7=> "000000000000000000000001000000010000000000000000000000000000000000000",  --Komentaro vieta
8=> "111010000010000000000000000000000000000000000000000000000000000000000",  --Komentaro vieta
9=> "000100000000000000000000000000000000000000000000000000000000000000000",  --Komentaro vieta
10=> "000000001000000000000000000000000000000000000000001000000000000000000",  --Komentaro vieta
11=> "001000000000000000000000000000000000000000000000000000000000000000000",  --Komentaro vieta
12=> "000000000000000100000000000000000000000000000000000000000000000000000",  --Komentaro vieta
13=> "000000100000000000000000000000000000000000000000000000000000000000000",  --Komentaro vieta
14=> "000000001000000000000000000000000000000000000000000001000000000000000",  --Komentaro vieta
15=> "001000000000000000000000000000000000000000000000000000000000000000000",  --Komentaro vieta
16=> "000000000000000000000010000000000000000000000000000000000000000000000",  --Komentaro vieta
17=> "000000100000000000000000000000000000000000000000000000000000000000000",  --Komentaro vieta
18=> "000000001000000000000000000000000000000000000000000100000000000000000",  --Komentaro vieta
19=> "001000000000000000000000000000000000000000000000000000000000000000000",  --Komentaro vieta
20=> "000000000000000000000000000000000000100000000000000000000000000000000",  --Komentaro vieta
21=> "010000000000000000000000000000000000000000010000000000000000000000000",  --Komentaro vieta
22=> "000000000000000000000001000000000000010000001000000000000000000000000",  --Komentaro vieta
23=> "000000000000000000000001000000000000010000001000000000000000000000000",  --Komentaro vieta
24=> "000000000000000000000001000000000000010000001000000000000000000000000",  --Komentaro vieta
25=> "000000000000000000000001000000000000010000001000000000000000000000000",  --Komentaro vieta
26=> "000000000000000000000001000000000000010000001000000000000000000000000",  --Komentaro vieta
27=> "000000000000000000000001000000000000010000001000000000000000000000000",  --Komentaro vieta
28=> "000000000000000000000001000000000000010000001000000000000000000000000",  --Komentaro vieta
29=> "000000000000000000000000000000000000000000001000000000000000000000000",  --Komentaro vieta
30=> "000100000000000000000000000000000000000000000000000000000010000000000",  --Komentaro vieta
31=> "000000001000000000000000000000000000000000000000001000000000000000000",  --Komentaro vieta
32=> "000010000000000000000000000000000000000000000000000000000000000010000",  --Komentaro vieta
33=> "000010001000000000000000000000000000000000000000001000000000000000000",  --Komentaro vieta
34=> "000000100000000000000000000000000000000000000000000000000000000000000",  --Komentaro vieta
35=> "100010010011100000000000000000000000000000000000000000000000000000000",  --Komentaro vieta
36=> "000000101000000000000000000000000000000000001000001000000000000000000",  --Komentaro vieta
37=> "000010000000000000000000000000000000000000000000000000000000000000000",  --Komentaro vieta
38=> "111110010100100000000000000000000000000000000000000000000000000000000",  --Komentaro vieta
39=> "000000000000000000000000000000000000000000000000100000000000000000000",  --Komentaro vieta
40=> "111110010100100000000000000000000000000000000000000000000000000000000",  --Komentaro vieta
41=> "000000000000000000000000000000000000000000000000000000000000000000001",  --Komentaro vieta
42=> "000000000100000000000000000000000000000000000000000000000000000000000",  --Komentaro vieta
43=> "111010010000100000000000000000000000000000000000000000000000000000000",  --Komentaro vieta
44=> "000000010000000000000000000000000000000000000000000000000000000000000",  --Komentaro vieta
45=> "000000001000000000000000000000000000000000000000000000100000000000000",  --Komentaro vieta
46=> "000000000000000000000000000000000000000000000000000000000000000000010",  --Komentaro vieta





	
	others => (others => '0') );   
	
	
	
begin
	process (RST_ROM, clk) 
		
	begin
		if RST_ROM'event and RST_ROM = '1' then 
			ROM_Dout <= ROM_CMDln(0);
		elsif clk'event and clk = '0' then
			ROM_Dout <= ROM_CMDln(to_integer(unsigned(ROM_CMD))); 
		end if;
		
	end process;
	
end rtl;